//MultMod
module MultTest
(input         clk , 
 input         rstn, 
 input         start,

 input[255:0]  aa    ,
 input[255:0]  bb    ,
 output[255:0] d
 );


reg[15:0] A[15:0],B[15:0],T[31:0],M[31:0],DD[15:0],MM[15:0],M3[31:0],TM[15:0],MT1,MT0,MT14,MT15,TT15;

reg[15:0] h0[15:0],l0[15:0],h1[15:0],l1[15:0],h2[15:0],l2[15:0],h3[15:0],l3[15:0],h4[15:0],l4[15:0],h5[15:0],l5[15:0],h6[15:0],l6[15:0],h7[15:0],l7[15:0],h8[15:0],l8[15:0],h9[15:0],l9[15:0],h10[15:0],l10[15:0],h11[15:0],l11[15:0],h12[15:0],l12[15:0],h13[15:0],l13[15:0],h14[15:0],l14[15:0],h15[15:0],l15[15:0];

reg[3:0] MT[16:0]; 
reg[4:0] T3[31:0];

reg[15:0]inv16,inv17,inv18,inv19,inv26,inv27,inv28,inv29,invT16,invT17,invT18,invT19,invT26,invT27,invT28,invT29;
reg[5:0]i;
reg[255:0] out; 
reg[261:0] out1,out2,out3;

reg[15:0] Asave, Bsave;
always@(posedge clk)
if(!rstn)
begin
    Asave<=16'h1234;
    Bsave<=16'h1234;
end
else
begin
    Asave<=aa[15:0];
    Bsave<=bb[15:0];
end

reg[15:0] Bsel0, Bsel1, Bsel2, Bsel3;
//test
parameter zero=16'h0000;

reg[1:0] clkNum, clkNum2;

//`ifdef DEBUG
wire[511:0] T3w, M3w;
assign T3w= {T3[31],T3[30],T3[29],T3[28],T3[27],T3[26],T3[25],T3[24],T3[23],T3[22],T3[21],T3[20],T3[19],T3[18],T3[17],T3[16],T3[15],T3[14],T3[13],T3[12],T3[11],T3[10],T3[9],T3[8],T3[7],T3[6],T3[5],T3[4],T3[3],T3[2],T3[1],T3[0]};
assign M3w= {M3[31],M3[30],M3[29],M3[28],M3[27],M3[26],M3[25],M3[24],M3[23],M3[22],M3[21],M3[20],M3[19],M3[18],M3[17],M3[16],M3[15],M3[14],M3[13],M3[12],M3[11],M3[10],M3[9],M3[8],M3[7],M3[6],M3[5],M3[4],M3[3],M3[2],M3[1],M3[0]};
//`endif

//assign Num=clkNum;
//reg [1:0]state,nextstate;
//parameter idle=2'd0,busy=2'd1;
reg flag_new;
always@(posedge clk)
if(!rstn)
    flag_new<=0;
else if((bb[15:0]!=Bsave) || (aa[15:0]!=Asave))
    flag_new<=1;
else 
    flag_new<=0;

reg flag_end;
always@(posedge clk)
    flag_end<=(clkNum==0);

always@(posedge clk)
  begin
    if(!rstn)// ||(!start))
      clkNum2<=4'b0;
    else if((bb[15:0]!=Bsave) || (aa[15:0]!=Asave))
      clkNum2<=4'b1;
    else if(clkNum2!=0)
      clkNum2<=clkNum2+4'b1;
  end

always@(posedge clk)
    clkNum<=clkNum2;
//cycle 1
always@(*)
begin
    A[0] =aa[15:0];
    A[1] =aa[31:16];
    A[2] =aa[47:32];
    A[3] =aa[63:48];
    A[4] =aa[79:64];
    A[5] =aa[95:80];
    A[6] =aa[111:96];
    A[7] =aa[127:112];
    A[8] =aa[143:128];
    A[9] =aa[159:144];
    A[10]=aa[175:160];
    A[11]=aa[191:176];
    A[12]=aa[207:192];
    A[13]=aa[223:208];
    A[14]=aa[239:224];
    A[15]=aa[255:240];
    
    B[0] =bb[15:0];
    B[1] =bb[31:16];
    B[2] =bb[47:32];
    B[3] =bb[63:48];
    B[4] =bb[79:64];
    B[5] =bb[95:80];
    B[6] =bb[111:96];
    B[7] =bb[127:112];
    B[8] =bb[143:128];
    B[9] =bb[159:144];
    B[10]=bb[175:160];
    B[11]=bb[191:176];
    B[12]=bb[207:192];
    B[13]=bb[223:208];
    B[14]=bb[239:224];
    B[15]=bb[255:240];
end

//cycle 2
always@(posedge clk)
for(i=0;i<16;i=i+1)
begin
    {h0[i],l0[i]}<=A[i]*B[0];
    {h1[i],l1[i]}<=A[i]*B[1];
    {h2[i],l2[i]}<=A[i]*B[2];
    {h3[i],l3[i]}<=A[i]*B[3];
    {h4[i],l4[i]}<=A[i]*B[4];
    {h5[i],l5[i]}<=A[i]*B[5];
    {h6[i],l6[i]}<=A[i]*B[6];
    {h7[i],l7[i]}<=A[i]*B[7];
    {h8[i],l8[i]}<=A[i]*B[8];
    {h9[i],l9[i]}<=A[i]*B[9];
    {h10[i],l10[i]}<=A[i]*B[10];
    {h11[i],l11[i]}<=A[i]*B[11];
    {h12[i],l12[i]}<=A[i]*B[12];
    {h13[i],l13[i]}<=A[i]*B[13];
    {h14[i],l14[i]}<=A[i]*B[14];
    {h15[i],l15[i]}<=A[i]*B[15];
end


wire[20:0] Tw0,Tw1,Tw2,Tw3,Tw4,Tw5,Tw6,Tw7,Tw8,Tw9,Tw10,Tw11,Tw12,Tw13,Tw14,Tw15,Tw16,Tw17,Tw18,Tw19,Tw20,Tw21,Tw22,Tw23,Tw24,Tw25,Tw26,Tw27,Tw28,Tw29,Tw30,Tw31;

assign Tw0=l0[0];
assign Tw2=l0[2]+l1[1]+h0[1]+l2[0]+h1[0];
assign Tw3=l0[3]+l1[2]+h0[2]+l2[1]+h1[1]+l3[0]+h2[0];
assign Tw4=l0[4]+l1[3]+h0[3]+l2[2]+h1[2]+l3[1]+h2[1]+l4[0]+h3[0];
assign Tw5=l0[5]+l1[4]+h0[4]+l2[3]+h1[3]+l3[2]+h2[2]+l4[1]+h3[1]+l5[0]+h4[0];
assign Tw6=l0[6]+l1[5]+h0[5]+l2[4]+h1[4]+l3[3]+h2[3]+l4[2]+h3[2]+l5[1]+h4[1]+l6[0]+h5[0];
assign Tw7=l0[7]+l1[6]+h0[6]+l2[5]+h1[5]+l3[4]+h2[4]+l4[3]+h3[3]+l5[2]+h4[2]+l6[1]+h5[1]+l7[0]+h6[0];
assign Tw8=l0[8]+l1[7]+h0[7]+l2[6]+h1[6]+l3[5]+h2[5]+l4[4]+h3[4]+l5[3]+h4[3]+l6[2]+h5[2]+l7[1]+h6[1]+l8[0]+h7[0];
assign Tw9=l0[9]+l1[8]+h0[8]+l2[7]+h1[7]+l3[6]+h2[6]+l4[5]+h3[5]+l5[4]+h4[4]+l6[3]+h5[3]+l7[2]+h6[2]+l8[1]+h7[1]+l9[0]+h8[0];
assign Tw10=l0[10]+l1[9]+h0[9]+l2[8]+h1[8]+l3[7]+h2[7]+l4[6]+h3[6]+l5[5]+h4[5]+l6[4]+h5[4]+l7[3]+h6[3]+l8[2]+h7[2]+l9[1]+h8[1]+l10[0]+h9[0];
assign Tw11=l0[11]+l1[10]+h0[10]+l2[9]+h1[9]+l3[8]+h2[8]+l4[7]+h3[7]+l5[6]+h4[6]+l6[5]+h5[5]+l7[4]+h6[4]+l8[3]+h7[3]+l9[2]+h8[2]+l10[1]+h9[1]+l11[0]+h10[0];
assign Tw12=l0[12]+l1[11]+h0[11]+l2[10]+h1[10]+l3[9]+h2[9]+l4[8]+h3[8]+l5[7]+h4[7]+l6[6]+h5[6]+l7[5]+h6[5]+l8[4]+h7[4]+l9[3]+h8[3]+l10[2]+h9[2]+l11[1]+h10[1]+l12[0]+h11[0];
assign Tw13=l0[13]+l1[12]+h0[12]+l2[11]+h1[11]+l3[10]+h2[10]+l4[9]+h3[9]+l5[8]+h4[8]+l6[7]+h5[7]+l7[6]+h6[6]+l8[5]+h7[5]+l9[4]+h8[4]+l10[3]+h9[3]+l11[2]+h10[2]+l12[1]+h11[1]+l13[0]+h12[0];
assign Tw14=l0[14]+l1[13]+h0[13]+l2[12]+h1[12]+l3[11]+h2[11]+l4[10]+h3[10]+l5[9]+h4[9]+l6[8]+h5[8]+l7[7]+h6[7]+l8[6]+h7[6]+l9[5]+h8[5]+l10[4]+h9[4]+l11[3]+h10[3]+l12[2]+h11[2]+l13[1]+h12[1]+l14[0]+h13[0];
assign Tw15=l0[15]+l1[14]+h0[14]+l2[13]+h1[13]+l3[12]+h2[12]+l4[11]+h3[11]+l5[10]+h4[10]+l6[9]+h5[9]+l7[8]+h6[8]+l8[7]+h7[7]+l9[6]+h8[6]+l10[5]+h9[5]+l11[4]+h10[4]+l12[3]+h11[3]+l13[2]+h12[2]+l14[1]+h13[1]+l15[0]+h14[0];
assign Tw16=l1[15]+h0[15]+l2[14]+h1[14]+l3[13]+h2[13]+l4[12]+h3[12]+l5[11]+h4[11]+l6[10]+h5[10]+l7[9]+h6[9]+l8[8]+h7[8]+l9[7]+h8[7]+l10[6]+h9[6]+l11[5]+h10[5]+l12[4]+h11[4]+l13[3]+h12[3]+l14[2]+h13[2]+l15[1]+h14[1]+h15[0];
assign Tw17=l2[15]+h1[15]+l3[14]+h2[14]+l4[13]+h3[13]+l5[12]+h4[12]+l6[11]+h5[11]+l7[10]+h6[10]+l8[9]+h7[9]+l9[8]+h8[8]+l10[7]+h9[7]+l11[6]+h10[6]+l12[5]+h11[5]+l13[4]+h12[4]+l14[3]+h13[3]+l15[2]+h14[2]+h15[1];
assign Tw18=l3[15]+h2[15]+l4[14]+h3[14]+l5[13]+h4[13]+l6[12]+h5[12]+l7[11]+h6[11]+l8[10]+h7[10]+l9[9]+h8[9]+l10[8]+h9[8]+l11[7]+h10[7]+l12[6]+h11[6]+l13[5]+h12[5]+l14[4]+h13[4]+l15[3]+h14[3]+h15[2];
assign Tw19=l4[15]+h3[15]+l5[14]+h4[14]+l6[13]+h5[13]+l7[12]+h6[12]+l8[11]+h7[11]+l9[10]+h8[10]+l10[9]+h9[9]+l11[8]+h10[8]+l12[7]+h11[7]+l13[6]+h12[6]+l14[5]+h13[5]+l15[4]+h14[4]+h15[3];
assign Tw20=l5[15]+h4[15]+l6[14]+h5[14]+l7[13]+h6[13]+l8[12]+h7[12]+l9[11]+h8[11]+l10[10]+h9[10]+l11[9]+h10[9]+l12[8]+h11[8]+l13[7]+h12[7]+l14[6]+h13[6]+l15[5]+h14[5]+h15[4];
assign Tw21=l6[15]+h5[15]+l7[14]+h6[14]+l8[13]+h7[13]+l9[12]+h8[12]+l10[11]+h9[11]+l11[10]+h10[10]+l12[9]+h11[9]+l13[8]+h12[8]+l14[7]+h13[7]+l15[6]+h14[6]+h15[5];
assign Tw22=l7[15]+h6[15]+l8[14]+h7[14]+l9[13]+h8[13]+l10[12]+h9[12]+l11[11]+h10[11]+l12[10]+h11[10]+l13[9]+h12[9]+l14[8]+h13[8]+l15[7]+h14[7]+h15[6];
assign Tw23=l8[15]+h7[15]+l9[14]+h8[14]+l10[13]+h9[13]+l11[12]+h10[12]+l12[11]+h11[11]+l13[10]+h12[10]+l14[9]+h13[9]+l15[8]+h14[8]+h15[7];
assign Tw24=l9[15]+h8[15]+l10[14]+h9[14]+l11[13]+h10[13]+l12[12]+h11[12]+l13[11]+h12[11]+l14[10]+h13[10]+l15[9]+h14[9]+h15[8];
assign Tw25=l10[15]+h9[15]+l11[14]+h10[14]+l12[13]+h11[13]+l13[12]+h12[12]+l14[11]+h13[11]+l15[10]+h14[10]+h15[9];
assign Tw26=l11[15]+h10[15]+l12[14]+h11[14]+l13[13]+h12[13]+l14[12]+h13[12]+l15[11]+h14[11]+h15[10];
assign Tw27=l12[15]+h11[15]+l13[14]+h12[14]+l14[13]+h13[13]+l15[12]+h14[12]+h15[11];
assign Tw28=l13[15]+h12[15]+l14[14]+h13[14]+l15[13]+h14[13]+h15[12];
assign Tw29=l14[15]+h13[15]+l15[14]+h14[14]+h15[13];
assign Tw30=l15[15]+h14[15]+h15[14];
assign Tw31=h15[15];


always @(posedge clk) 
begin
    {T3[0],M3[0]}<=Tw0;
    {T3[1],M3[1]}<=Tw1;
    {T3[2],M3[2]}<=Tw2;
    {T3[3],M3[3]}<=Tw3;
    {T3[4],M3[4]}<=Tw4;
    {T3[5],M3[5]}<=Tw5;
    {T3[6],M3[6]}<=Tw6;
    {T3[7],M3[7]}<=Tw7;
    {T3[8],M3[8]}<=Tw8;
    {T3[9],M3[9]}<=Tw9;
    {T3[11],M3[11]}<=Tw11;
    {T3[12],M3[12]}<=Tw12;
    {T3[13],M3[13]}<=Tw13;
    {T3[14],M3[14]}<=Tw14;
    {T3[15],M3[15]}<=Tw15;
    {T3[16],M3[16]}<=Tw16;
    {T3[17],M3[17]}<=Tw17;
    {T3[18],M3[18]}<=Tw18;
    {T3[19],M3[19]}<=Tw19;
    {T3[20],M3[20]}<=Tw20;
    {T3[21],M3[21]}<=Tw21;
    {T3[22],M3[22]}<=Tw22;
    {T3[23],M3[23]}<=Tw23;
    {T3[24],M3[24]}<=Tw24;
    {T3[25],M3[25]}<=Tw25;
    {T3[26],M3[26]}<=Tw26;
    {T3[27],M3[27]}<=Tw27;
    {T3[28],M3[28]}<=Tw28;
    {T3[29],M3[29]}<=Tw29;
    {T3[30],M3[30]}<=Tw30;
    {T3[31],M3[31]}<=Tw31;
end

//cycle 5
always@(*)  
begin
    inv16=~M3[16];inv17=~M3[17];inv18=~M3[18];inv19=~M3[19];inv26=~M3[26];inv27=~M3[27];inv28=~M3[28];inv29=~M3[29];
    invT16=~T3[15];invT17=~T3[16];invT18=~T3[17];invT19=~T3[18];invT26=~T3[25];invT27=~T3[26];invT28=~T3[27];invT29=~T3[28];  
end

always@(posedge clk)
//if(flag_end)
begin
    {MT[0],MM[0]}<=M3[0]+{M3[26],1'b0}+{M3[30],1'b0}+{M3[28],1'b0}+M3[16]+M3[18]+M3[22]+M3[24]+M3[20]+
    {T3[25],1'b0}+{T3[29],1'b0}+{T3[27],1'b0}+T3[15]+T3[17]+T3[21]+T3[23]+T3[19];

    {MT[1],MM[1]}<=M3[1]+{M3[27],1'b0}+{M3[31],1'b0}+{M3[29],1'b0}+M3[17]+M3[19]+M3[23]+M3[25]+M3[21] +
    T3[0]+{T3[26],1'b0}+{T3[30],1'b0}+{T3[28],1'b0}+T3[16]+T3[18]+T3[22]+T3[24]+T3[20];

    {MT[2],MM[2]}<=M3[2]+M3[28]+M3[30]+M3[28]+M3[30]+M3[26]+M3[18]+M3[20]+M3[22]+M3[24]+
    T3[1]+T3[27]+T3[29]+T3[27]+T3[29]+T3[25]+T3[17]+T3[19]+T3[21]+T3[23];

    {MT[3],MM[3]}<=M3[3]+M3[29]+M3[31]+M3[29]+M3[31]+M3[27]+M3[19]+M3[23]+M3[25]+M3[21]+
    T3[2]+T3[28]+T3[30]+T3[28]+T3[30]+T3[26]+T3[18]+T3[22]+T3[24]+T3[20];

    {MT[4],MM[4]}<=M3[4]+16'd4+inv16+inv18+inv26+inv28+
    T3[3]+16'h4+invT16+invT18+invT26+invT28;

    {MT[5],MM[5]}<=M3[5]+inv17+inv19+inv27+inv29+
    T3[4]+invT17+invT19+invT27+invT29;

    {MT[6],MM[6]}<=M3[6]+M3[26]+M3[26]+M3[22]+M3[24]+M3[28]+M3[30]+M3[16]+16'hfffc+
    T3[5]+{T3[25],1'b0}+T3[21]+T3[23]+T3[27]+T3[29]+T3[15]+16'hfffc;

    {MT[7],MM[7]}<=M3[7]+M3[27]+M3[27]+M3[23]+M3[25]+M3[29]+M3[31]+M3[17]+16'hffff+
    T3[6]+T3[26]+T3[26]+T3[22]+T3[24]+T3[28]+T3[30]+T3[16]+16'hffff;

    {MT[8],MM[8]}<=M3[8]+M3[28]+M3[28]+M3[30]+M3[26]+M3[18]+M3[24]+16'hffff+
    T3[7]+T3[27]+T3[27]+T3[29]+T3[25]+T3[17]+T3[23]+16'hffff;

    {MT[9],MM[9]}<=M3[9]+M3[29]+M3[29]+M3[31]+M3[27]+M3[19]+M3[25]+16'hffff+
    T3[8]+T3[28]+T3[28]+T3[30]+T3[26]+T3[18]+T3[24]+16'hffff;

    {MT[10],MM[10]}<=M3[10]+M3[30]+M3[30]+M3[28]+M3[26]+M3[20]+16'hffff+
    T3[9]+T3[29]+T3[29]+T3[27]+T3[25]+T3[19]+16'hffff;

    {MT[11],MM[11]}<=M3[11]+M3[31]+M3[31]+M3[29]+M3[27]+M3[21]+16'hffff+
    T3[10]+T3[30]+T3[30]+T3[28]+T3[26]+T3[20]+16'hffff;

    {MT[12],MM[12]}<=M3[12]+M3[30]+M3[28]+M3[22]+16'hffff+
    T3[11]+T3[29]+T3[27]+T3[21]+16'hffff;

    {MT[13],MM[13]}<=M3[13]+M3[31]+M3[29]+M3[23]+16'hffff+
    T3[12]+T3[30]+T3[28]+T3[22]+16'hffff;

    {MT[14],MM[14]}<=M3[14]+M3[16]+M3[18]+M3[20]+M3[22]+{M3[24],1'b0}+{M3[26],1'b0}+{M3[28],1'b0}+{M3[30],1'b0}+M3[30]+16'hffff+
                    T3[13]+T3[15]+T3[17]+T3[19]+T3[21]+{T3[23],1'b0}+{T3[25],1'b0}+{T3[27],1'b0}+{T3[29],1'b0}+T3[29]+16'hffff;

    {MT[15],MM[15]}<=M3[15]+M3[17]+M3[19]+M3[21]+M3[23]+{M3[25],1'b0}+{M3[27],1'b0}+{M3[29],1'b0}+{M3[31],1'b0}+M3[31]+16'hffff+
                    T3[14]+T3[16]+T3[18]+T3[20]+T3[22]+{T3[24],1'b0}+{T3[26],1'b0}+{T3[28],1'b0}+{T3[30],1'b0}+T3[30]+16'hffff;
end   

reg cor; //correction bit, in case that out1[127:0] exceeds 128-bit
//cycle 6
always@(*)   
begin
    out1[261:128] = {17'h1fffe,MM[15],MM[14],MM[13],MM[12],MM[11],MM[10],MM[9],MM[8]}+
            {MT[15],12'h0, MT[14],12'h0, MT[13],12'h0, MT[12],12'h0, MT[11],12'h0, MT[10],12'h0, MT[9],12'h0, MT[8], 12'h0, MT[7]};
    
    {cor, out1[127:0]} = {MM[7],MM[6],MM[5],MM[4],MM[3],MM[2],MM[1],MM[0]}+
            {MT[6],12'h0, MT[5],12'h0, MT[4],12'h0, MT[3],12'h0, MT[2],12'h0, MT[1],12'h0, MT[0], 16'h0};
              
end

reg[5:0] out2_hi, out2_hi2;
always@(posedge clk)    
begin
    out2[261:0]<=out1[261:0];  
    out2_hi<=(out1[128+15: 128]==16'hffff)? out1[261:256]+cor : out1[261:256];
    out2_hi2<= (out1[128+15: 128]==16'hffff)? cor :0;
end 

//cycle 7  
always@(posedge clk) 
begin
    out[63:0] <= out2[63:0]+ out2_hi;
    out[255-32:64] <= out2[255-32:64] - out2_hi +{out2_hi, 32'h0}+{out2_hi2, 64'b0};
    out[255: 255-31] <= out2[255: 255-31] + out2_hi + out2_hi2;
end
 
assign d=out[255:0];

endmodule